package isa_decls_bh(
    package isa_defines
    ,package isa_decls_bh
) where

import isa_defines

type XLEN_2 = TMul XLEN 2
type XLEN_MINUS_2 = TSub XLEN 2

xlen:: Integer
xlen = valueOf XLEN

data RVVersion = RV32 | RV64 deriving (Eq, Bits)
rv_version:: RVVersion
rv_version = case xlen of {
    32 -> RV32;
    64 -> RV64;
}

type BitsPerByte = 8
type Byte = Bit BitsPerByte
bits_per_byte:: Integer
bits_per_byte = valueOf BitsPerByte

type BitsPerWordXL = XLEN
type WordXL = Bit BitsPerWordXL

type BytesPerWordXL = TDiv BitsPerWordXL BitsPerByte
bytes_per_wordxl:: Integer
bytes_per_wordxl = valueOf BytesPerWordXL

type Bits_per_Byte_in_WordXL = TLog BytesPerWordXL
type Byte_in_WordXL = Bit Bits_per_Byte_in_WordXL
bits_per_byte_in_wordxl:: Integer
bits_per_byte_in_wordxl = valueOf Bits_per_Byte_in_WordXL

type IntXL = Int XLEN
type Addr = WordXL

{-
// ================================================================
// FLEN and related constants, for floating point data
// Can have one or two fpu sizes (should they be merged sooner than later ?).

// ISA_D => ISA_F (ISA_D implies ISA_F)
// The combination ISA_D and !ISA_F is not permitted
-}

type WordFL = Bit FLEN
type BytesPerWordFL = TDiv FLEN BitsPerByte

{-
// ================================================================
// Tokens are used for signalling/synchronization, and have no payload
-}
type Token = Bit 0

{-
// ================================================================
// Instruction fields
// This is used for encoding Tandem Verifier traces
-}
data ISize = ISIZE16 | ISIZE32 deriving (Bits, Eq, FShow)

type InstrBits = Bit 32
type Opcode = Bit 7
type RegIdx = Bit 5
type CSRAddr = Bit 12

type NumRegs = 32
num_regs:: Integer
num_regs = valueOf NumRegs

illegal_instr:: InstrBits
illegal_instr = 32'h0000_0000

instr_opcode:: InstrBits -> Opcode
instr_opcode x = x[6:0]

instr_funct2:: InstrBits -> Bit 2
instr_funct2 x = x[26:25]
instr_funct3:: InstrBits -> Bit 3
instr_funct3 x = x[14:12]
instr_funct5:: InstrBits -> Bit 5
instr_funct5 x = x[31:27]
instr_funct7:: InstrBits -> Bit 7
instr_funct7 x = x[31:25]
instr_funct10:: InstrBits -> Bit 10
instr_funct10 x = x[31:25] ++ x[14:12]
instr_fmt:: InstrBits -> Bit 2
instr_fmt x = x[26:25]

instr_rd:: InstrBits -> RegIdx
instr_rd x = x[11:7]
instr_rs1:: InstrBits -> RegIdx
instr_rs1 x = x[19:15]
instr_rs2:: InstrBits -> RegIdx
instr_rs2 x = x[24:20]
instr_rs3:: InstrBits -> RegIdx
instr_rs3 x =  x[31:27]
instr_csr:: InstrBits -> CSRAddr
instr_csr x = x[31:20]
instr_I_imm12:: InstrBits -> Bit 12
instr_I_imm12 x = x[31:20]
instr_S_imm12:: InstrBits -> Bit 12
instr_S_imm12 x = x[31:25] ++ x[11:7]
instr_U_imm20:: InstrBits -> Bit 20
instr_U_imm20 x = x[31:12]

instr_B_imm13:: InstrBits -> Bit 13
instr_B_imm13 x = x[31:31] ++ x[7:7] ++ x[30:25] ++ x[11:8] ++ 1'b0

instr_J_imm21:: InstrBits -> Bit 21
instr_J_imm21 x = x[31:31] ++ x[19:12] ++ x [20:20] ++ x[30:21] ++ 1'b0

-- For FENCE decode
instr_pred:: InstrBits -> Bit 4
instr_pred x = x[27:24]
instr_succ:: InstrBits -> Bit 4
instr_succ x = x[23:20]

-- For AMO decode
instr_aqrl:: InstrBits -> Bit 2
instr_aqrl x = x[26:25]

data InstrFmt = InstrFmtNone | InstrFmtR | InstrFmtI 
    deriving (Bits, Eq, FShow)

-- difference with haskell, semicolon ; is used to seperation
data InstrType = Raw InstrBits | R {
    funct7:: (Bit 7);
    rs2:: RegIdx;
    rs1:: RegIdx;
    funct3:: Bit 3;
    rd:: RegIdx;
    opcode:: Opcode;
} | I {
    imm12:: Bit 12;
    rs1:: RegIdx;
    funct3:: Bit 3;
    rd:: RegIdx;
    opcode:: Opcode;
} deriving (Bits, FShow)

-- difference with haskell, `struct` keyword is used for record type instead of data
struct Instruction = {
    fmt:: InstrFmt;
    ast:: InstrType;
} deriving (Bits, FShow)

decode_instruction:: InstrBits -> Instruction
decode_instruction x = case x[6:0] of {
    7'b0110011 -> Instruction {fmt = InstrFmtR; ast = R (unpack x)};
    7'b0010011 -> Instruction {fmt = InstrFmtI; ast = I (unpack x)};
    _ -> Instruction {fmt = InstrFmtNone; ast = Raw x};
}

encode_instr_R:: Bit 7 -> RegIdx -> RegIdx -> Bit 3 -> RegIdx -> Bit 7 -> InstrBits
encode_instr_R funct7 rs2 rs1 funct3 rd opcode = 
    funct7 ++ rs2 ++ rs1 ++ funct3 ++ rd ++ opcode

encode_instr_I:: Bit 12 -> RegIdx -> Bit 3 -> RegIdx -> Opcode -> InstrBits
encode_instr_I imm12 rs1 funct3 rd opcode = 
    imm12 ++ rs1 ++ funct3 ++ rd ++ opcode

encode_instr_S:: Bit 12 -> RegIdx -> RegIdx -> Bit 3 -> Opcode -> InstrBits
encode_instr_S imm12 rs2 rs1 funct3 opcode = 
    imm12[11:5] ++ rs2 ++ rs1 ++ funct3 ++ imm12[4:0] ++ opcode

encode_instr_B:: Bit 13 -> RegIdx -> RegIdx -> Bit 3 -> Opcode -> InstrBits
encode_instr_B imm13 rs2 rs1 funct3 opcode = 
    imm13[12:12] ++ imm13[10:5] ++ rs2 ++ rs1 ++ funct3 ++ imm13[4:1] ++ imm13[11:11] ++ opcode

encode_instr_U:: Bit 20 -> RegIdx -> Opcode -> InstrBits
encode_instr_U imm20 rd opcode = imm20 ++ rd ++ opcode

encode_instr_J:: Bit 21 -> RegIdx -> Opcode -> InstrBits
encode_instr_J imm21 rd opcode = 
    imm21[20:20] ++ imm21[10:1] ++ imm21[11:11] ++ imm21[19:12] ++ rd ++ opcode
