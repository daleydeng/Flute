package defines_bh;
#include "defines.bsvi"
endpackage