package GPR_RegFile(
   GPR_RegFile_IFC (..) 
   ,mkGPR_RegFile) where

import RegFile
import ClientServer
import FIFOF
import GetPut
import GetPut_Aux

import isa_types

interface GPR_RegFile_IFC =
   server_reset:: Server Token Token

   read_rs1:: RegIdx -> WordXL
   read_rs1_port2:: RegIdx -> WordXL -- For debugger access only
   read_rs2:: RegIdx -> WordXL 
   write_rd:: RegIdx -> WordXL -> Action

data RF_State = RF_RESET_START | RF_RESETTING | RF_RUNNING deriving (Eq, Bits, FShow);

mkGPR_RegFile:: Module GPR_RegFile_IFC
mkGPR_RegFile = 
   module
      rg_state:: Reg RF_State <- mkReg RF_RESET_START
      f_reset_rsps:: FIFOF Token <- mkFIFOF

      -- General Purpose Registers
      -- TODO: can we use Reg [0] for some other purpose?
      regfile::RegFile RegIdx WordXL <- mkRegFileFull

--    -- ----------------------------------------------------------------
--    -- Reset.
--    -- This loop initializes all GPRs to 0.
--    -- The spec does not require this, but it's useful for debugging
--    -- and tandem verification

-- `ifdef INCLUDE_TANDEM_VERIF
      rg_j:: Reg RegIdx <- mkRegU    -- reset loop index
-- #endif

      rules
         "rl_reset_start": when rg_state == RF_RESET_START
            ==> action rg_state := RF_RESETTING

         "rl_reset_loop": when rg_state == RF_RESETTING, kINCLUDE_TANDEM_VERIF == 0
            ==> action rg_state := RF_RUNNING

         "rl_reset_start": when rg_state == RF_RESET_START, kINCLUDE_TANDEM_VERIF == 1
            ==> action rg_j := 1

         "rl_reset_loop": when rg_state == RF_RESETTING, kINCLUDE_TANDEM_VERIF == 1
            ==> action
                  regfile.upd rg_j 0;
                  rg_j := rg_j + 1;
                  case rg_j of 31 -> rg_state := RF_RUNNING 


      mk_server_reset_request:: Put Token
      mk_server_reset_request <- 
         module 
            interface
               put token = action 
                  rg_state := RF_RESET_START
                  -- This response is placed here, and not in rl_reset_loop, because
                  -- reset_loop can happen on power-up, where no response is expected.
                  f_reset_rsps.enq token

      mk_server_reset_response:: Get Token
      mk_server_reset_response <- 
         module
            interface
               get = pop f_reset_rsps when rg_state == RF_RUNNING

      mk_server_reset:: Server Token Token
      mk_server_reset <-
         module 
            interface
               request = mk_server_reset_request
               response = mk_server_reset_response

      interface
         server_reset = mk_server_reset
         server_reset = mk_server_reset

         read_rs1 rs1 = if rs1 == 0 then 0 else regfile.sub rs1

         read_rs1_port2 rs1 = if rs1 == 0 then 0 else regfile.sub rs1
         read_rs2 rs2 = if rs2 == 0 then 0 else regfile.sub rs2
         write_rd rd rd_val = rd != 0 ?? regfile.upd rd rd_val when rg_state == RF_RUNNING
