// Copyright (c) 2016-2022 Bluespec, Inc. All Rights Reserved

package CPU_IFC;

// ================================================================
// BSV library imports

import GetPut       :: *;
import ClientServer :: *;

// ================================================================
// Project imports

import isa_base :: *;

import AXI4_Types   :: *;
import AXI_Widths   :: *;    // For Wd_Id/Addr/Data/User_Dma
import Fabric_Defs  :: *;
import Near_Mem_IFC :: *;

#ifdef INCLUDE_DMEM_SLAVE
import AXI4_Lite_Types :: *;
#endif

#ifdef INCLUDE_GDB_CONTROL
import DM_CPU_Req_Rsp :: *;
#endif

#ifdef INCLUDE_PC_TRACE
import PCTrace :: *;
#endif

#ifdef INCLUDE_TANDEM_VERIF
import tv_trace_data :: *;
#endif

// ================================================================
// CPU interface

interface CPU_IFC;
   // Reset
   interface Server #(Bool, Bool)  hart0_server_reset;

   // ----------------
   // SoC fabric connections

   // IMem to Fabric master interface
   interface AXI4_Master_IFC #(Wd_Id, Wd_Addr, Wd_Data, Wd_User)  imem_master;

   // Fabric master interface to memory
   interface Near_Mem_Fabric_IFC  mem_master;

   // ----------------------------------------------------------------
   // Optional AXI4-Lite D-cache slave interface

#ifdef INCLUDE_DMEM_SLAVE
   interface AXI4_Lite_Slave_IFC #(Wd_Addr, Wd_Data, Wd_User)  dmem_slave;
#endif

   // ----------------
   // Interface to 'coherent DMA' port of optional L2 cache

   interface AXI4_Slave_IFC #(Wd_Id_Dma, Wd_Addr_Dma, Wd_Data_Dma, Wd_User_Dma)  dma_server;

   // ----------------------------------------------------------------
   // External interrupts

   (* always_ready, always_enabled *)
   method Action  m_external_interrupt_req (Bool set_not_clear);

   (* always_ready, always_enabled *)
   method Action  s_external_interrupt_req (Bool set_not_clear);

   // ----------------
   // Set CSR TIME (shadow-copy of MTIME)

   (* always_ready, always_enabled *)
   method Action ma_set_csr_time (Bit#(64) t);

   // ----------------
   // Software and timer interrupts (from Near_Mem_IO/CLINT)

   (* always_ready, always_enabled *)
   method Action  software_interrupt_req (Bool set_not_clear);

   (* always_ready, always_enabled *)
   method Action  timer_interrupt_req    (Bool set_not_clear);

   // ----------------
   // Non-maskable interrupt

   (* always_ready, always_enabled *)
   method Action  nmi_req (Bool set_not_clear);

   // ----------------
   // Optional PC trace interface
   // Outputs a stream of 2-tuples: (cycle_count, pc)

#ifdef INCLUDE_PC_TRACE
   interface Get #(PCTrace)  g_pc_trace;
#endif

   // ----------------
   // Optional interface to Tandem Verifier

#ifdef INCLUDE_TANDEM_VERIF
   interface Get #(TraceData)  trace_data_out;
#endif

   // ----------------
   // Optional interface to Debug Module

#ifdef INCLUDE_GDB_CONTROL
   // run-control, other
   interface Server #(Bool, Bool)  hart0_server_run_halt;
   interface Put #(Bit#(4))       hart0_put_other_req;

   // GPR access
   interface Server #(DM_CPU_Req #(5,  XLEN), DM_CPU_Rsp #(XLEN)) hart0_gpr_mem_server;

#ifdef ISA_F
   // FPR access
   interface Server #(DM_CPU_Req #(5,  FLEN), DM_CPU_Rsp #(FLEN)) hart0_fpr_mem_server;
#endif

   // CSR access
   interface Server #(DM_CPU_Req #(12, XLEN), DM_CPU_Rsp #(XLEN)) hart0_csr_mem_server;
#endif

   // ----------------------------------------------------------------
   // Misc. control and status

   // ----------------
   // Debugging: set core's verbosity

   method Action set_verbosity (Bit#(4)  verbosity, Bit#(64)  logdelay);

   // ----------------
   // For ISA tests: watch memory writes to <tohost> addr

#ifdef WATCH_TOHOST
   method Action set_watch_tohost (Bool watch_tohost, Bit#(64) tohost_addr);
   method Bit#(64) mv_tohost_value;
#endif

   // Inform core that DDR4 has been initialized and is ready to accept requests
   method Action ma_ddr4_ready;

   // Misc. status; 0 = running, no error
   (* always_ready *)
   method Bit#(8) mv_status;

endinterface

// ================================================================

endpackage
