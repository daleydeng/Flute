package isa_defines_bh;
`include "isa_defines.bsvi"
endpackage