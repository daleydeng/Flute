package isa_defines;

`include "isa_defines.bsvi"

endpackage